`timescale 1ns/1ps

module twiddle_tb();

endmodule 